`ifndef RES_NET_PKG
`define RES_NET_PKG

package RES_NET_PKG;

// Codebook_C = [[-1,  1, -1, -1, -1, -1,  1, -1, -1, -1,  1,  1,  1, -1, -1,  1, -1,  1, -1,  1,  1, -1, -1, -1, -1, -1, -1,  1, -1,  1, -1,  1],
//               [ 1, -1, -1,  1,  1, -1, -1, -1, -1,  1,  1,  1,  1, -1,  1, -1, -1, -1,  1,  1, -1, -1,  1,  1,  1, -1,  1,  1, -1, -1, -1,  1],
//               [ 1,  1,  1,  1, -1, -1,  1,  1,  1, -1,  1,  1, -1,  1, -1,  1, -1,  1,  1, -1, -1,  1, -1,  1,  1, -1,  1,  1,  1, -1, -1,  1]]   
parameter VECTOR_LEN = 32;
parameter NUM_CODEBOOK_BITS = 4;
// Color Codebook times its transpose
parameter logic signed [VECTOR_LEN-1 : 0][VECTOR_LEN-1 : 0][NUM_CODEBOOK_BITS-1 : 0] CCT = {{4'b0011, 4'b1111, 4'b0001, 4'b0001, 4'b0001, 4'b1101, 4'b0011, 4'b0001, 4'b1101, 4'b0001, 4'b1111, 4'b0001, 4'b0001, 4'b0001, 4'b1101, 4'b1111, 4'b1111, 4'b1101, 4'b0001, 4'b0001, 4'b0001, 4'b0001, 4'b0001, 4'b0001, 4'b0011, 4'b0001, 4'b1111, 4'b1101, 4'b1111, 4'b1111, 4'b1101, 4'b0001},
                                                                               {4'b1111, 4'b0011, 4'b0001, 4'b0001, 4'b0001, 4'b0001, 4'b1111, 4'b1101, 4'b0001, 4'b0001, 4'b0011, 4'b0001, 4'b1101, 4'b0001, 4'b0001, 4'b1111, 4'b1111, 4'b0001, 4'b1101, 4'b1101, 4'b1101, 4'b1101, 4'b0001, 4'b1101, 4'b1111, 4'b0001, 4'b0011, 4'b0001, 4'b0011, 4'b1111, 4'b0001, 4'b0001},
                                                                               {4'b0001, 4'b0001, 4'b0011, 4'b1111, 4'b1111, 4'b1111, 4'b0001, 4'b1111, 4'b1111, 4'b1111, 4'b0001, 4'b0011, 4'b1111, 4'b1111, 4'b1111, 4'b0001, 4'b0001, 4'b1111, 4'b1111, 4'b1111, 4'b1111, 4'b1111, 4'b0011, 4'b1111, 4'b0001, 4'b1111, 4'b0001, 4'b1111, 4'b0001, 4'b0001, 4'b1111, 4'b0011},
                                                                               {4'b0001, 4'b0001, 4'b1111, 4'b0011, 4'b0011, 4'b1111, 4'b0001, 4'b1111, 4'b1111, 4'b0011, 4'b0001, 4'b1111, 4'b1111, 4'b0011, 4'b1111, 4'b1101, 4'b1101, 4'b1111, 4'b1111, 4'b1111, 4'b1111, 4'b1111, 4'b1111, 4'b1111, 4'b0001, 4'b0011, 4'b0001, 4'b1111, 4'b0001, 4'b1101, 4'b1111, 4'b1111},
                                                                               {4'b0001, 4'b0001, 4'b1111, 4'b0011, 4'b0011, 4'b1111, 4'b0001, 4'b1111, 4'b1111, 4'b0011, 4'b0001, 4'b1111, 4'b1111, 4'b0011, 4'b1111, 4'b1101, 4'b1101, 4'b1111, 4'b1111, 4'b1111, 4'b1111, 4'b1111, 4'b1111, 4'b1111, 4'b0001, 4'b0011, 4'b0001, 4'b1111, 4'b0001, 4'b1101, 4'b1111, 4'b1111},
                                                                               {4'b1101, 4'b0001, 4'b1111, 4'b1111, 4'b1111, 4'b0011, 4'b1101, 4'b1111, 4'b0011, 4'b1111, 4'b0001, 4'b1111, 4'b1111, 4'b1111, 4'b0011, 4'b0001, 4'b0001, 4'b0011, 4'b1111, 4'b1111, 4'b1111, 4'b1111, 4'b1111, 4'b1111, 4'b1101, 4'b1111, 4'b0001, 4'b0011, 4'b0001, 4'b0001, 4'b0011, 4'b1111},
                                                                               {4'b0011, 4'b1111, 4'b0001, 4'b0001, 4'b0001, 4'b1101, 4'b0011, 4'b0001, 4'b1101, 4'b0001, 4'b1111, 4'b0001, 4'b0001, 4'b0001, 4'b1101, 4'b1111, 4'b1111, 4'b1101, 4'b0001, 4'b0001, 4'b0001, 4'b0001, 4'b0001, 4'b0001, 4'b0011, 4'b0001, 4'b1111, 4'b1101, 4'b1111, 4'b1111, 4'b1101, 4'b0001},
                                                                               {4'b0001, 4'b1101, 4'b1111, 4'b1111, 4'b1111, 4'b1111, 4'b0001, 4'b0011, 4'b1111, 4'b1111, 4'b1101, 4'b1111, 4'b0011, 4'b1111, 4'b1111, 4'b0001, 4'b0001, 4'b1111, 4'b0011, 4'b0011, 4'b0011, 4'b0011, 4'b1111, 4'b0011, 4'b0001, 4'b1111, 4'b1101, 4'b1111, 4'b1101, 4'b0001, 4'b1111, 4'b1111},
                                                                               {4'b1101, 4'b0001, 4'b1111, 4'b1111, 4'b1111, 4'b0011, 4'b1101, 4'b1111, 4'b0011, 4'b1111, 4'b0001, 4'b1111, 4'b1111, 4'b1111, 4'b0011, 4'b0001, 4'b0001, 4'b0011, 4'b1111, 4'b1111, 4'b1111, 4'b1111, 4'b1111, 4'b1111, 4'b1101, 4'b1111, 4'b0001, 4'b0011, 4'b0001, 4'b0001, 4'b0011, 4'b1111},
                                                                               {4'b0001, 4'b0001, 4'b1111, 4'b0011, 4'b0011, 4'b1111, 4'b0001, 4'b1111, 4'b1111, 4'b0011, 4'b0001, 4'b1111, 4'b1111, 4'b0011, 4'b1111, 4'b1101, 4'b1101, 4'b1111, 4'b1111, 4'b1111, 4'b1111, 4'b1111, 4'b1111, 4'b1111, 4'b0001, 4'b0011, 4'b0001, 4'b1111, 4'b0001, 4'b1101, 4'b1111, 4'b1111},
                                                                               {4'b1111, 4'b0011, 4'b0001, 4'b0001, 4'b0001, 4'b0001, 4'b1111, 4'b1101, 4'b0001, 4'b0001, 4'b0011, 4'b0001, 4'b1101, 4'b0001, 4'b0001, 4'b1111, 4'b1111, 4'b0001, 4'b1101, 4'b1101, 4'b1101, 4'b1101, 4'b0001, 4'b1101, 4'b1111, 4'b0001, 4'b0011, 4'b0001, 4'b0011, 4'b1111, 4'b0001, 4'b0001},
                                                                               {4'b0001, 4'b0001, 4'b0011, 4'b1111, 4'b1111, 4'b1111, 4'b0001, 4'b1111, 4'b1111, 4'b1111, 4'b0001, 4'b0011, 4'b1111, 4'b1111, 4'b1111, 4'b0001, 4'b0001, 4'b1111, 4'b1111, 4'b1111, 4'b1111, 4'b1111, 4'b0011, 4'b1111, 4'b0001, 4'b1111, 4'b0001, 4'b1111, 4'b0001, 4'b0001, 4'b1111, 4'b0011},
                                                                               {4'b0001, 4'b1101, 4'b1111, 4'b1111, 4'b1111, 4'b1111, 4'b0001, 4'b0011, 4'b1111, 4'b1111, 4'b1101, 4'b1111, 4'b0011, 4'b1111, 4'b1111, 4'b0001, 4'b0001, 4'b1111, 4'b0011, 4'b0011, 4'b0011, 4'b0011, 4'b1111, 4'b0011, 4'b0001, 4'b1111, 4'b1101, 4'b1111, 4'b1101, 4'b0001, 4'b1111, 4'b1111},
                                                                               {4'b0001, 4'b0001, 4'b1111, 4'b0011, 4'b0011, 4'b1111, 4'b0001, 4'b1111, 4'b1111, 4'b0011, 4'b0001, 4'b1111, 4'b1111, 4'b0011, 4'b1111, 4'b1101, 4'b1101, 4'b1111, 4'b1111, 4'b1111, 4'b1111, 4'b1111, 4'b1111, 4'b1111, 4'b0001, 4'b0011, 4'b0001, 4'b1111, 4'b0001, 4'b1101, 4'b1111, 4'b1111},
                                                                               {4'b1101, 4'b0001, 4'b1111, 4'b1111, 4'b1111, 4'b0011, 4'b1101, 4'b1111, 4'b0011, 4'b1111, 4'b0001, 4'b1111, 4'b1111, 4'b1111, 4'b0011, 4'b0001, 4'b0001, 4'b0011, 4'b1111, 4'b1111, 4'b1111, 4'b1111, 4'b1111, 4'b1111, 4'b1101, 4'b1111, 4'b0001, 4'b0011, 4'b0001, 4'b0001, 4'b0011, 4'b1111},
                                                                               {4'b1111, 4'b1111, 4'b0001, 4'b1101, 4'b1101, 4'b0001, 4'b1111, 4'b0001, 4'b0001, 4'b1101, 4'b1111, 4'b0001, 4'b0001, 4'b1101, 4'b0001, 4'b0011, 4'b0011, 4'b0001, 4'b0001, 4'b0001, 4'b0001, 4'b0001, 4'b0001, 4'b0001, 4'b1111, 4'b1101, 4'b1111, 4'b0001, 4'b1111, 4'b0011, 4'b0001, 4'b0001},
                                                                               {4'b1111, 4'b1111, 4'b0001, 4'b1101, 4'b1101, 4'b0001, 4'b1111, 4'b0001, 4'b0001, 4'b1101, 4'b1111, 4'b0001, 4'b0001, 4'b1101, 4'b0001, 4'b0011, 4'b0011, 4'b0001, 4'b0001, 4'b0001, 4'b0001, 4'b0001, 4'b0001, 4'b0001, 4'b1111, 4'b1101, 4'b1111, 4'b0001, 4'b1111, 4'b0011, 4'b0001, 4'b0001},
                                                                               {4'b1101, 4'b0001, 4'b1111, 4'b1111, 4'b1111, 4'b0011, 4'b1101, 4'b1111, 4'b0011, 4'b1111, 4'b0001, 4'b1111, 4'b1111, 4'b1111, 4'b0011, 4'b0001, 4'b0001, 4'b0011, 4'b1111, 4'b1111, 4'b1111, 4'b1111, 4'b1111, 4'b1111, 4'b1101, 4'b1111, 4'b0001, 4'b0011, 4'b0001, 4'b0001, 4'b0011, 4'b1111},
                                                                               {4'b0001, 4'b1101, 4'b1111, 4'b1111, 4'b1111, 4'b1111, 4'b0001, 4'b0011, 4'b1111, 4'b1111, 4'b1101, 4'b1111, 4'b0011, 4'b1111, 4'b1111, 4'b0001, 4'b0001, 4'b1111, 4'b0011, 4'b0011, 4'b0011, 4'b0011, 4'b1111, 4'b0011, 4'b0001, 4'b1111, 4'b1101, 4'b1111, 4'b1101, 4'b0001, 4'b1111, 4'b1111},
                                                                               {4'b0001, 4'b1101, 4'b1111, 4'b1111, 4'b1111, 4'b1111, 4'b0001, 4'b0011, 4'b1111, 4'b1111, 4'b1101, 4'b1111, 4'b0011, 4'b1111, 4'b1111, 4'b0001, 4'b0001, 4'b1111, 4'b0011, 4'b0011, 4'b0011, 4'b0011, 4'b1111, 4'b0011, 4'b0001, 4'b1111, 4'b1101, 4'b1111, 4'b1101, 4'b0001, 4'b1111, 4'b1111},
                                                                               {4'b0001, 4'b1101, 4'b1111, 4'b1111, 4'b1111, 4'b1111, 4'b0001, 4'b0011, 4'b1111, 4'b1111, 4'b1101, 4'b1111, 4'b0011, 4'b1111, 4'b1111, 4'b0001, 4'b0001, 4'b1111, 4'b0011, 4'b0011, 4'b0011, 4'b0011, 4'b1111, 4'b0011, 4'b0001, 4'b1111, 4'b1101, 4'b1111, 4'b1101, 4'b0001, 4'b1111, 4'b1111},
                                                                               {4'b0001, 4'b1101, 4'b1111, 4'b1111, 4'b1111, 4'b1111, 4'b0001, 4'b0011, 4'b1111, 4'b1111, 4'b1101, 4'b1111, 4'b0011, 4'b1111, 4'b1111, 4'b0001, 4'b0001, 4'b1111, 4'b0011, 4'b0011, 4'b0011, 4'b0011, 4'b1111, 4'b0011, 4'b0001, 4'b1111, 4'b1101, 4'b1111, 4'b1101, 4'b0001, 4'b1111, 4'b1111},
                                                                               {4'b0001, 4'b0001, 4'b0011, 4'b1111, 4'b1111, 4'b1111, 4'b0001, 4'b1111, 4'b1111, 4'b1111, 4'b0001, 4'b0011, 4'b1111, 4'b1111, 4'b1111, 4'b0001, 4'b0001, 4'b1111, 4'b1111, 4'b1111, 4'b1111, 4'b1111, 4'b0011, 4'b1111, 4'b0001, 4'b1111, 4'b0001, 4'b1111, 4'b0001, 4'b0001, 4'b1111, 4'b0011},
                                                                               {4'b0001, 4'b1101, 4'b1111, 4'b1111, 4'b1111, 4'b1111, 4'b0001, 4'b0011, 4'b1111, 4'b1111, 4'b1101, 4'b1111, 4'b0011, 4'b1111, 4'b1111, 4'b0001, 4'b0001, 4'b1111, 4'b0011, 4'b0011, 4'b0011, 4'b0011, 4'b1111, 4'b0011, 4'b0001, 4'b1111, 4'b1101, 4'b1111, 4'b1101, 4'b0001, 4'b1111, 4'b1111},
                                                                               {4'b0011, 4'b1111, 4'b0001, 4'b0001, 4'b0001, 4'b1101, 4'b0011, 4'b0001, 4'b1101, 4'b0001, 4'b1111, 4'b0001, 4'b0001, 4'b0001, 4'b1101, 4'b1111, 4'b1111, 4'b1101, 4'b0001, 4'b0001, 4'b0001, 4'b0001, 4'b0001, 4'b0001, 4'b0011, 4'b0001, 4'b1111, 4'b1101, 4'b1111, 4'b1111, 4'b1101, 4'b0001},
                                                                               {4'b0001, 4'b0001, 4'b1111, 4'b0011, 4'b0011, 4'b1111, 4'b0001, 4'b1111, 4'b1111, 4'b0011, 4'b0001, 4'b1111, 4'b1111, 4'b0011, 4'b1111, 4'b1101, 4'b1101, 4'b1111, 4'b1111, 4'b1111, 4'b1111, 4'b1111, 4'b1111, 4'b1111, 4'b0001, 4'b0011, 4'b0001, 4'b1111, 4'b0001, 4'b1101, 4'b1111, 4'b1111},
                                                                               {4'b1111, 4'b0011, 4'b0001, 4'b0001, 4'b0001, 4'b0001, 4'b1111, 4'b1101, 4'b0001, 4'b0001, 4'b0011, 4'b0001, 4'b1101, 4'b0001, 4'b0001, 4'b1111, 4'b1111, 4'b0001, 4'b1101, 4'b1101, 4'b1101, 4'b1101, 4'b0001, 4'b1101, 4'b1111, 4'b0001, 4'b0011, 4'b0001, 4'b0011, 4'b1111, 4'b0001, 4'b0001},
                                                                               {4'b1101, 4'b0001, 4'b1111, 4'b1111, 4'b1111, 4'b0011, 4'b1101, 4'b1111, 4'b0011, 4'b1111, 4'b0001, 4'b1111, 4'b1111, 4'b1111, 4'b0011, 4'b0001, 4'b0001, 4'b0011, 4'b1111, 4'b1111, 4'b1111, 4'b1111, 4'b1111, 4'b1111, 4'b1101, 4'b1111, 4'b0001, 4'b0011, 4'b0001, 4'b0001, 4'b0011, 4'b1111},
                                                                               {4'b1111, 4'b0011, 4'b0001, 4'b0001, 4'b0001, 4'b0001, 4'b1111, 4'b1101, 4'b0001, 4'b0001, 4'b0011, 4'b0001, 4'b1101, 4'b0001, 4'b0001, 4'b1111, 4'b1111, 4'b0001, 4'b1101, 4'b1101, 4'b1101, 4'b1101, 4'b0001, 4'b1101, 4'b1111, 4'b0001, 4'b0011, 4'b0001, 4'b0011, 4'b1111, 4'b0001, 4'b0001},
                                                                               {4'b1111, 4'b1111, 4'b0001, 4'b1101, 4'b1101, 4'b0001, 4'b1111, 4'b0001, 4'b0001, 4'b1101, 4'b1111, 4'b0001, 4'b0001, 4'b1101, 4'b0001, 4'b0011, 4'b0011, 4'b0001, 4'b0001, 4'b0001, 4'b0001, 4'b0001, 4'b0001, 4'b0001, 4'b1111, 4'b1101, 4'b1111, 4'b0001, 4'b1111, 4'b0011, 4'b0001, 4'b0001},
                                                                               {4'b1101, 4'b0001, 4'b1111, 4'b1111, 4'b1111, 4'b0011, 4'b1101, 4'b1111, 4'b0011, 4'b1111, 4'b0001, 4'b1111, 4'b1111, 4'b1111, 4'b0011, 4'b0001, 4'b0001, 4'b0011, 4'b1111, 4'b1111, 4'b1111, 4'b1111, 4'b1111, 4'b1111, 4'b1101, 4'b1111, 4'b0001, 4'b0011, 4'b0001, 4'b0001, 4'b0011, 4'b1111},
                                                                               {4'b0001, 4'b0001, 4'b0011, 4'b1111, 4'b1111, 4'b1111, 4'b0001, 4'b1111, 4'b1111, 4'b1111, 4'b0001, 4'b0011, 4'b1111, 4'b1111, 4'b1111, 4'b0001, 4'b0001, 4'b1111, 4'b1111, 4'b1111, 4'b1111, 4'b1111, 4'b0011, 4'b1111, 4'b0001, 4'b1111, 4'b0001, 4'b1111, 4'b0001, 4'b0001, 4'b1111, 4'b0011}};


// Codebook_S = [[-1, -1,  1,  1,  1, -1, -1,  1,  1,  1, -1, -1,  1,  1, -1,  1, -1, -1,  1, -1,  1, -1, -1, -1, -1, -1, -1,  1, -1, -1,  1,  1],
//               [ 1,  1,  1,  1,  1, -1, -1,  1,  1, -1,  1, -1, -1, -1,  1, -1, -1, -1, -1,  1,  1, -1, -1, -1,  1, -1, -1, -1,  1,  1, -1, -1],
//               [-1,  1, -1, -1,  1,  1,  1, -1,  1,  1,  1,  1, -1,  1,  1, -1, -1, -1,  1, -1, -1, -1, -1, -1, -1, -1,  1,  1,  1,  1,  1, -1]]

// Shape Codebook times its transpose
parameter logic signed [VECTOR_LEN-1 : 0][VECTOR_LEN-1 : 0][NUM_CODEBOOK_BITS-1 : 0] SST = {{4'b0011, 4'b1111, 4'b1111, 4'b0001, 4'b0001, 4'b0011, 4'b0011, 4'b1111, 4'b0001, 4'b0001, 4'b0011, 4'b0001, 4'b1111, 4'b0001, 4'b0001, 4'b0011, 4'b0001, 4'b1111, 4'b1101, 4'b0001, 4'b0001, 4'b1111, 4'b0011, 4'b1111, 4'b0001, 4'b1111, 4'b1101, 4'b1101, 4'b0001, 4'b1111, 4'b0001, 4'b0001},
                                                                                            {4'b1111, 4'b0011, 4'b1111, 4'b1101, 4'b1101, 4'b1111, 4'b1111, 4'b1111, 4'b1101, 4'b0001, 4'b1111, 4'b0001, 4'b1111, 4'b1101, 4'b0001, 4'b1111, 4'b0001, 4'b0011, 4'b0001, 4'b0001, 4'b1101, 4'b0011, 4'b1111, 4'b0011, 4'b0001, 4'b1111, 4'b0001, 4'b0001, 4'b1101, 4'b0011, 4'b0001, 4'b1101},
                                                                                            {4'b1111, 4'b1111, 4'b0011, 4'b0001, 4'b0001, 4'b1111, 4'b1111, 4'b1111, 4'b0001, 4'b1101, 4'b1111, 4'b0001, 4'b0011, 4'b0001, 4'b0001, 4'b1111, 4'b1101, 4'b1111, 4'b0001, 4'b0001, 4'b0001, 4'b1111, 4'b1111, 4'b1111, 4'b0001, 4'b1111, 4'b0001, 4'b0001, 4'b0001, 4'b1111, 4'b0001, 4'b0001},
                                                                                            {4'b0001, 4'b1101, 4'b0001, 4'b0011, 4'b0011, 4'b0001, 4'b0001, 4'b0001, 4'b0011, 4'b1111, 4'b0001, 4'b1111, 4'b0001, 4'b0011, 4'b1111, 4'b0001, 4'b1111, 4'b1101, 4'b1111, 4'b1111, 4'b0011, 4'b1101, 4'b0001, 4'b1101, 4'b1111, 4'b0001, 4'b1111, 4'b1111, 4'b0011, 4'b1101, 4'b1111, 4'b0011},
                                                                                            {4'b0001, 4'b1101, 4'b0001, 4'b0011, 4'b0011, 4'b0001, 4'b0001, 4'b0001, 4'b0011, 4'b1111, 4'b0001, 4'b1111, 4'b0001, 4'b0011, 4'b1111, 4'b0001, 4'b1111, 4'b1101, 4'b1111, 4'b1111, 4'b0011, 4'b1101, 4'b0001, 4'b1101, 4'b1111, 4'b0001, 4'b1111, 4'b1111, 4'b0011, 4'b1101, 4'b1111, 4'b0011},
                                                                                            {4'b0011, 4'b1111, 4'b1111, 4'b0001, 4'b0001, 4'b0011, 4'b0011, 4'b1111, 4'b0001, 4'b0001, 4'b0011, 4'b0001, 4'b1111, 4'b0001, 4'b0001, 4'b0011, 4'b0001, 4'b1111, 4'b1101, 4'b0001, 4'b0001, 4'b1111, 4'b0011, 4'b1111, 4'b0001, 4'b1111, 4'b1101, 4'b1101, 4'b0001, 4'b1111, 4'b0001, 4'b0001},
                                                                                            {4'b0011, 4'b1111, 4'b1111, 4'b0001, 4'b0001, 4'b0011, 4'b0011, 4'b1111, 4'b0001, 4'b0001, 4'b0011, 4'b0001, 4'b1111, 4'b0001, 4'b0001, 4'b0011, 4'b0001, 4'b1111, 4'b1101, 4'b0001, 4'b0001, 4'b1111, 4'b0011, 4'b1111, 4'b0001, 4'b1111, 4'b1101, 4'b1101, 4'b0001, 4'b1111, 4'b0001, 4'b0001},
                                                                                            {4'b1111, 4'b1111, 4'b1111, 4'b0001, 4'b0001, 4'b1111, 4'b1111, 4'b0011, 4'b0001, 4'b0001, 4'b1111, 4'b1101, 4'b1111, 4'b0001, 4'b1101, 4'b1111, 4'b0001, 4'b1111, 4'b0001, 4'b1101, 4'b0001, 4'b1111, 4'b1111, 4'b1111, 4'b1101, 4'b0011, 4'b0001, 4'b0001, 4'b0001, 4'b1111, 4'b1101, 4'b0001},
                                                                                            {4'b0001, 4'b1101, 4'b0001, 4'b0011, 4'b0011, 4'b0001, 4'b0001, 4'b0001, 4'b0011, 4'b1111, 4'b0001, 4'b1111, 4'b0001, 4'b0011, 4'b1111, 4'b0001, 4'b1111, 4'b1101, 4'b1111, 4'b1111, 4'b0011, 4'b1101, 4'b0001, 4'b1101, 4'b1111, 4'b0001, 4'b1111, 4'b1111, 4'b0011, 4'b1101, 4'b1111, 4'b0011},
                                                                                            {4'b0001, 4'b0001, 4'b1101, 4'b1111, 4'b1111, 4'b0001, 4'b0001, 4'b0001, 4'b1111, 4'b0011, 4'b0001, 4'b1111, 4'b1101, 4'b1111, 4'b1111, 4'b0001, 4'b0011, 4'b0001, 4'b1111, 4'b1111, 4'b1111, 4'b0001, 4'b0001, 4'b0001, 4'b1111, 4'b0001, 4'b1111, 4'b1111, 4'b1111, 4'b0001, 4'b1111, 4'b1111},
                                                                                            {4'b0011, 4'b1111, 4'b1111, 4'b0001, 4'b0001, 4'b0011, 4'b0011, 4'b1111, 4'b0001, 4'b0001, 4'b0011, 4'b0001, 4'b1111, 4'b0001, 4'b0001, 4'b0011, 4'b0001, 4'b1111, 4'b1101, 4'b0001, 4'b0001, 4'b1111, 4'b0011, 4'b1111, 4'b0001, 4'b1111, 4'b1101, 4'b1101, 4'b0001, 4'b1111, 4'b0001, 4'b0001},
                                                                                            {4'b0001, 4'b0001, 4'b0001, 4'b1111, 4'b1111, 4'b0001, 4'b0001, 4'b1101, 4'b1111, 4'b1111, 4'b0001, 4'b0011, 4'b0001, 4'b1111, 4'b0011, 4'b0001, 4'b1111, 4'b0001, 4'b1111, 4'b0011, 4'b1111, 4'b0001, 4'b0001, 4'b0001, 4'b0011, 4'b1101, 4'b1111, 4'b1111, 4'b1111, 4'b0001, 4'b0011, 4'b1111},
                                                                                            {4'b1111, 4'b1111, 4'b0011, 4'b0001, 4'b0001, 4'b1111, 4'b1111, 4'b1111, 4'b0001, 4'b1101, 4'b1111, 4'b0001, 4'b0011, 4'b0001, 4'b0001, 4'b1111, 4'b1101, 4'b1111, 4'b0001, 4'b0001, 4'b0001, 4'b1111, 4'b1111, 4'b1111, 4'b0001, 4'b1111, 4'b0001, 4'b0001, 4'b0001, 4'b1111, 4'b0001, 4'b0001},
                                                                                            {4'b0001, 4'b1101, 4'b0001, 4'b0011, 4'b0011, 4'b0001, 4'b0001, 4'b0001, 4'b0011, 4'b1111, 4'b0001, 4'b1111, 4'b0001, 4'b0011, 4'b1111, 4'b0001, 4'b1111, 4'b1101, 4'b1111, 4'b1111, 4'b0011, 4'b1101, 4'b0001, 4'b1101, 4'b1111, 4'b0001, 4'b1111, 4'b1111, 4'b0011, 4'b1101, 4'b1111, 4'b0011},
                                                                                            {4'b0001, 4'b0001, 4'b0001, 4'b1111, 4'b1111, 4'b0001, 4'b0001, 4'b1101, 4'b1111, 4'b1111, 4'b0001, 4'b0011, 4'b0001, 4'b1111, 4'b0011, 4'b0001, 4'b1111, 4'b0001, 4'b1111, 4'b0011, 4'b1111, 4'b0001, 4'b0001, 4'b0001, 4'b0011, 4'b1101, 4'b1111, 4'b1111, 4'b1111, 4'b0001, 4'b0011, 4'b1111},
                                                                                            {4'b0011, 4'b1111, 4'b1111, 4'b0001, 4'b0001, 4'b0011, 4'b0011, 4'b1111, 4'b0001, 4'b0001, 4'b0011, 4'b0001, 4'b1111, 4'b0001, 4'b0001, 4'b0011, 4'b0001, 4'b1111, 4'b1101, 4'b0001, 4'b0001, 4'b1111, 4'b0011, 4'b1111, 4'b0001, 4'b1111, 4'b1101, 4'b1101, 4'b0001, 4'b1111, 4'b0001, 4'b0001},
                                                                                            {4'b0001, 4'b0001, 4'b1101, 4'b1111, 4'b1111, 4'b0001, 4'b0001, 4'b0001, 4'b1111, 4'b0011, 4'b0001, 4'b1111, 4'b1101, 4'b1111, 4'b1111, 4'b0001, 4'b0011, 4'b0001, 4'b1111, 4'b1111, 4'b1111, 4'b0001, 4'b0001, 4'b0001, 4'b1111, 4'b0001, 4'b1111, 4'b1111, 4'b1111, 4'b0001, 4'b1111, 4'b1111},
                                                                                            {4'b1111, 4'b0011, 4'b1111, 4'b1101, 4'b1101, 4'b1111, 4'b1111, 4'b1111, 4'b1101, 4'b0001, 4'b1111, 4'b0001, 4'b1111, 4'b1101, 4'b0001, 4'b1111, 4'b0001, 4'b0011, 4'b0001, 4'b0001, 4'b1101, 4'b0011, 4'b1111, 4'b0011, 4'b0001, 4'b1111, 4'b0001, 4'b0001, 4'b1101, 4'b0011, 4'b0001, 4'b1101},
                                                                                            {4'b1101, 4'b0001, 4'b0001, 4'b1111, 4'b1111, 4'b1101, 4'b1101, 4'b0001, 4'b1111, 4'b1111, 4'b1101, 4'b1111, 4'b0001, 4'b1111, 4'b1111, 4'b1101, 4'b1111, 4'b0001, 4'b0011, 4'b1111, 4'b1111, 4'b0001, 4'b1101, 4'b0001, 4'b1111, 4'b0001, 4'b0011, 4'b0011, 4'b1111, 4'b0001, 4'b1111, 4'b1111},
                                                                                            {4'b0001, 4'b0001, 4'b0001, 4'b1111, 4'b1111, 4'b0001, 4'b0001, 4'b1101, 4'b1111, 4'b1111, 4'b0001, 4'b0011, 4'b0001, 4'b1111, 4'b0011, 4'b0001, 4'b1111, 4'b0001, 4'b1111, 4'b0011, 4'b1111, 4'b0001, 4'b0001, 4'b0001, 4'b0011, 4'b1101, 4'b1111, 4'b1111, 4'b1111, 4'b0001, 4'b0011, 4'b1111},
                                                                                            {4'b0001, 4'b1101, 4'b0001, 4'b0011, 4'b0011, 4'b0001, 4'b0001, 4'b0001, 4'b0011, 4'b1111, 4'b0001, 4'b1111, 4'b0001, 4'b0011, 4'b1111, 4'b0001, 4'b1111, 4'b1101, 4'b1111, 4'b1111, 4'b0011, 4'b1101, 4'b0001, 4'b1101, 4'b1111, 4'b0001, 4'b1111, 4'b1111, 4'b0011, 4'b1101, 4'b1111, 4'b0011},
                                                                                            {4'b1111, 4'b0011, 4'b1111, 4'b1101, 4'b1101, 4'b1111, 4'b1111, 4'b1111, 4'b1101, 4'b0001, 4'b1111, 4'b0001, 4'b1111, 4'b1101, 4'b0001, 4'b1111, 4'b0001, 4'b0011, 4'b0001, 4'b0001, 4'b1101, 4'b0011, 4'b1111, 4'b0011, 4'b0001, 4'b1111, 4'b0001, 4'b0001, 4'b1101, 4'b0011, 4'b0001, 4'b1101},
                                                                                            {4'b0011, 4'b1111, 4'b1111, 4'b0001, 4'b0001, 4'b0011, 4'b0011, 4'b1111, 4'b0001, 4'b0001, 4'b0011, 4'b0001, 4'b1111, 4'b0001, 4'b0001, 4'b0011, 4'b0001, 4'b1111, 4'b1101, 4'b0001, 4'b0001, 4'b1111, 4'b0011, 4'b1111, 4'b0001, 4'b1111, 4'b1101, 4'b1101, 4'b0001, 4'b1111, 4'b0001, 4'b0001},
                                                                                            {4'b1111, 4'b0011, 4'b1111, 4'b1101, 4'b1101, 4'b1111, 4'b1111, 4'b1111, 4'b1101, 4'b0001, 4'b1111, 4'b0001, 4'b1111, 4'b1101, 4'b0001, 4'b1111, 4'b0001, 4'b0011, 4'b0001, 4'b0001, 4'b1101, 4'b0011, 4'b1111, 4'b0011, 4'b0001, 4'b1111, 4'b0001, 4'b0001, 4'b1101, 4'b0011, 4'b0001, 4'b1101},
                                                                                            {4'b0001, 4'b0001, 4'b0001, 4'b1111, 4'b1111, 4'b0001, 4'b0001, 4'b1101, 4'b1111, 4'b1111, 4'b0001, 4'b0011, 4'b0001, 4'b1111, 4'b0011, 4'b0001, 4'b1111, 4'b0001, 4'b1111, 4'b0011, 4'b1111, 4'b0001, 4'b0001, 4'b0001, 4'b0011, 4'b1101, 4'b1111, 4'b1111, 4'b1111, 4'b0001, 4'b0011, 4'b1111},
                                                                                            {4'b1111, 4'b1111, 4'b1111, 4'b0001, 4'b0001, 4'b1111, 4'b1111, 4'b0011, 4'b0001, 4'b0001, 4'b1111, 4'b1101, 4'b1111, 4'b0001, 4'b1101, 4'b1111, 4'b0001, 4'b1111, 4'b0001, 4'b1101, 4'b0001, 4'b1111, 4'b1111, 4'b1111, 4'b1101, 4'b0011, 4'b0001, 4'b0001, 4'b0001, 4'b1111, 4'b1101, 4'b0001},
                                                                                            {4'b1101, 4'b0001, 4'b0001, 4'b1111, 4'b1111, 4'b1101, 4'b1101, 4'b0001, 4'b1111, 4'b1111, 4'b1101, 4'b1111, 4'b0001, 4'b1111, 4'b1111, 4'b1101, 4'b1111, 4'b0001, 4'b0011, 4'b1111, 4'b1111, 4'b0001, 4'b1101, 4'b0001, 4'b1111, 4'b0001, 4'b0011, 4'b0011, 4'b1111, 4'b0001, 4'b1111, 4'b1111},
                                                                                            {4'b1101, 4'b0001, 4'b0001, 4'b1111, 4'b1111, 4'b1101, 4'b1101, 4'b0001, 4'b1111, 4'b1111, 4'b1101, 4'b1111, 4'b0001, 4'b1111, 4'b1111, 4'b1101, 4'b1111, 4'b0001, 4'b0011, 4'b1111, 4'b1111, 4'b0001, 4'b1101, 4'b0001, 4'b1111, 4'b0001, 4'b0011, 4'b0011, 4'b1111, 4'b0001, 4'b1111, 4'b1111},
                                                                                            {4'b0001, 4'b1101, 4'b0001, 4'b0011, 4'b0011, 4'b0001, 4'b0001, 4'b0001, 4'b0011, 4'b1111, 4'b0001, 4'b1111, 4'b0001, 4'b0011, 4'b1111, 4'b0001, 4'b1111, 4'b1101, 4'b1111, 4'b1111, 4'b0011, 4'b1101, 4'b0001, 4'b1101, 4'b1111, 4'b0001, 4'b1111, 4'b1111, 4'b0011, 4'b1101, 4'b1111, 4'b0011},
                                                                                            {4'b1111, 4'b0011, 4'b1111, 4'b1101, 4'b1101, 4'b1111, 4'b1111, 4'b1111, 4'b1101, 4'b0001, 4'b1111, 4'b0001, 4'b1111, 4'b1101, 4'b0001, 4'b1111, 4'b0001, 4'b0011, 4'b0001, 4'b0001, 4'b1101, 4'b0011, 4'b1111, 4'b0011, 4'b0001, 4'b1111, 4'b0001, 4'b0001, 4'b1101, 4'b0011, 4'b0001, 4'b1101},
                                                                                            {4'b0001, 4'b0001, 4'b0001, 4'b1111, 4'b1111, 4'b0001, 4'b0001, 4'b1101, 4'b1111, 4'b1111, 4'b0001, 4'b0011, 4'b0001, 4'b1111, 4'b0011, 4'b0001, 4'b1111, 4'b0001, 4'b1111, 4'b0011, 4'b1111, 4'b0001, 4'b0001, 4'b0001, 4'b0011, 4'b1101, 4'b1111, 4'b1111, 4'b1111, 4'b0001, 4'b0011, 4'b1111},
                                                                                            {4'b0001, 4'b1101, 4'b0001, 4'b0011, 4'b0011, 4'b0001, 4'b0001, 4'b0001, 4'b0011, 4'b1111, 4'b0001, 4'b1111, 4'b0001, 4'b0011, 4'b1111, 4'b0001, 4'b1111, 4'b1101, 4'b1111, 4'b1111, 4'b0011, 4'b1101, 4'b0001, 4'b1101, 4'b1111, 4'b0001, 4'b1111, 4'b1111, 4'b0011, 4'b1101, 4'b1111, 4'b0011}};




// Codebook_P = [[-1, -1,  1,  1, -1,  1, -1, -1, -1, -1,  1, -1, -1, -1, -1,  1, -1, -1,  1,  1, -1,  1,  1,  1, -1, -1, -1,  1,  1,  1,  1, -1],
//               [-1,  1, -1, -1,  1,  1, -1, -1, -1,  1, -1, -1, -1, -1, -1, -1, -1,  1,  1, -1,  1,  1, -1,  1,  1, -1, -1, -1,  1, -1, -1,  1],
//               [-1,  1, -1,  1,  1,  1, -1, -1,  1, -1,  1, -1,  1,  1,  1,  1,  1, -1, -1, -1, -1,  1, -1,  1,  1,  1, -1,  1, -1,  1, -1,  1],
//               [-1,  1,  1,  1,  1, -1, -1, -1, -1,  1,  1,  1,  1,  1, -1,  1,  1,  1,  1,  1,  1, -1, -1,  1,  1,  1,  1, -1,  1,  1,  1, -1]]

// Position Codebook times its transpose
parameter logic signed [VECTOR_LEN-1 : 0][VECTOR_LEN-1 : 0][NUM_CODEBOOK_BITS-1 : 0] PPT = {{4'b0100, 4'b0010, 4'b0010, 4'b0000, 4'b0010, 4'b0000, 4'b0100, 4'b0000, 4'b0000, 4'b0100, 4'b0000, 4'b0010, 4'b0000, 4'b1110, 4'b0010, 4'b0000, 4'b1110, 4'b1100, 4'b0010, 4'b0010, 4'b0010, 4'b1110, 4'b0000, 4'b1110, 4'b0000, 4'b0000, 4'b0100, 4'b0010, 4'b0000, 4'b1110, 4'b1100, 4'b0100},
                                                                                            {4'b0010, 4'b0100, 4'b0100, 4'b1110, 4'b0000, 4'b1110, 4'b0010, 4'b0010, 4'b0010, 4'b0010, 4'b1110, 4'b0000, 4'b1110, 4'b0000, 4'b0000, 4'b1110, 4'b0000, 4'b1110, 4'b0100, 4'b0000, 4'b0000, 4'b0000, 4'b0010, 4'b1100, 4'b1110, 4'b1110, 4'b0010, 4'b0000, 4'b1110, 4'b0000, 4'b1110, 4'b0010},
                                                                                            {4'b0010, 4'b0100, 4'b0100, 4'b1110, 4'b0000, 4'b1110, 4'b0010, 4'b0010, 4'b0010, 4'b0010, 4'b1110, 4'b0000, 4'b1110, 4'b0000, 4'b0000, 4'b1110, 4'b0000, 4'b1110, 4'b0100, 4'b0000, 4'b0000, 4'b0000, 4'b0010, 4'b1100, 4'b1110, 4'b1110, 4'b0010, 4'b0000, 4'b1110, 4'b0000, 4'b1110, 4'b0010},
                                                                                            {4'b0000, 4'b1110, 4'b1110, 4'b0100, 4'b0010, 4'b0100, 4'b0000, 4'b1100, 4'b1100, 4'b0000, 4'b0100, 4'b0010, 4'b0100, 4'b1110, 4'b0010, 4'b0100, 4'b1110, 4'b0000, 4'b1110, 4'b0010, 4'b0010, 4'b1110, 4'b0000, 4'b0010, 4'b0100, 4'b0000, 4'b0000, 4'b0010, 4'b0000, 4'b0010, 4'b0000, 4'b0000},
                                                                                            {4'b0010, 4'b0000, 4'b0000, 4'b0010, 4'b0100, 4'b0010, 4'b0010, 4'b1110, 4'b1110, 4'b0010, 4'b0010, 4'b0100, 4'b0010, 4'b1100, 4'b0100, 4'b0010, 4'b0000, 4'b1110, 4'b0000, 4'b0100, 4'b0100, 4'b1100, 4'b0010, 4'b0000, 4'b0010, 4'b0010, 4'b0010, 4'b0100, 4'b0010, 4'b0000, 4'b1110, 4'b0010},
                                                                                            {4'b0000, 4'b1110, 4'b1110, 4'b0100, 4'b0010, 4'b0100, 4'b0000, 4'b1100, 4'b1100, 4'b0000, 4'b0100, 4'b0010, 4'b0100, 4'b1110, 4'b0010, 4'b0100, 4'b1110, 4'b0000, 4'b1110, 4'b0010, 4'b0010, 4'b1110, 4'b0000, 4'b0010, 4'b0100, 4'b0000, 4'b0000, 4'b0010, 4'b0000, 4'b0010, 4'b0000, 4'b0000},
                                                                                            {4'b0100, 4'b0010, 4'b0010, 4'b0000, 4'b0010, 4'b0000, 4'b0100, 4'b0000, 4'b0000, 4'b0100, 4'b0000, 4'b0010, 4'b0000, 4'b1110, 4'b0010, 4'b0000, 4'b1110, 4'b1100, 4'b0010, 4'b0010, 4'b0010, 4'b1110, 4'b0000, 4'b1110, 4'b0000, 4'b0000, 4'b0100, 4'b0010, 4'b0000, 4'b1110, 4'b1100, 4'b0100},
                                                                                            {4'b0000, 4'b0010, 4'b0010, 4'b1100, 4'b1110, 4'b1100, 4'b0000, 4'b0100, 4'b0100, 4'b0000, 4'b1100, 4'b1110, 4'b1100, 4'b0010, 4'b1110, 4'b1100, 4'b0010, 4'b0000, 4'b0010, 4'b1110, 4'b1110, 4'b0010, 4'b0000, 4'b1110, 4'b1100, 4'b0000, 4'b0000, 4'b1110, 4'b0000, 4'b1110, 4'b0000, 4'b0000},
                                                                                            {4'b0000, 4'b0010, 4'b0010, 4'b1100, 4'b1110, 4'b1100, 4'b0000, 4'b0100, 4'b0100, 4'b0000, 4'b1100, 4'b1110, 4'b1100, 4'b0010, 4'b1110, 4'b1100, 4'b0010, 4'b0000, 4'b0010, 4'b1110, 4'b1110, 4'b0010, 4'b0000, 4'b1110, 4'b1100, 4'b0000, 4'b0000, 4'b1110, 4'b0000, 4'b1110, 4'b0000, 4'b0000},
                                                                                            {4'b0100, 4'b0010, 4'b0010, 4'b0000, 4'b0010, 4'b0000, 4'b0100, 4'b0000, 4'b0000, 4'b0100, 4'b0000, 4'b0010, 4'b0000, 4'b1110, 4'b0010, 4'b0000, 4'b1110, 4'b1100, 4'b0010, 4'b0010, 4'b0010, 4'b1110, 4'b0000, 4'b1110, 4'b0000, 4'b0000, 4'b0100, 4'b0010, 4'b0000, 4'b1110, 4'b1100, 4'b0100},
                                                                                            {4'b0000, 4'b1110, 4'b1110, 4'b0100, 4'b0010, 4'b0100, 4'b0000, 4'b1100, 4'b1100, 4'b0000, 4'b0100, 4'b0010, 4'b0100, 4'b1110, 4'b0010, 4'b0100, 4'b1110, 4'b0000, 4'b1110, 4'b0010, 4'b0010, 4'b1110, 4'b0000, 4'b0010, 4'b0100, 4'b0000, 4'b0000, 4'b0010, 4'b0000, 4'b0010, 4'b0000, 4'b0000},
                                                                                            {4'b0010, 4'b0000, 4'b0000, 4'b0010, 4'b0100, 4'b0010, 4'b0010, 4'b1110, 4'b1110, 4'b0010, 4'b0010, 4'b0100, 4'b0010, 4'b1100, 4'b0100, 4'b0010, 4'b0000, 4'b1110, 4'b0000, 4'b0100, 4'b0100, 4'b1100, 4'b0010, 4'b0000, 4'b0010, 4'b0010, 4'b0010, 4'b0100, 4'b0010, 4'b0000, 4'b1110, 4'b0010},
                                                                                            {4'b0000, 4'b1110, 4'b1110, 4'b0100, 4'b0010, 4'b0100, 4'b0000, 4'b1100, 4'b1100, 4'b0000, 4'b0100, 4'b0010, 4'b0100, 4'b1110, 4'b0010, 4'b0100, 4'b1110, 4'b0000, 4'b1110, 4'b0010, 4'b0010, 4'b1110, 4'b0000, 4'b0010, 4'b0100, 4'b0000, 4'b0000, 4'b0010, 4'b0000, 4'b0010, 4'b0000, 4'b0000},
                                                                                            {4'b1110, 4'b0000, 4'b0000, 4'b1110, 4'b1100, 4'b1110, 4'b1110, 4'b0010, 4'b0010, 4'b1110, 4'b1110, 4'b1100, 4'b1110, 4'b0100, 4'b1100, 4'b1110, 4'b0000, 4'b0010, 4'b0000, 4'b1100, 4'b1100, 4'b0100, 4'b1110, 4'b0000, 4'b1110, 4'b1110, 4'b1110, 4'b1100, 4'b1110, 4'b0000, 4'b0010, 4'b1110},
                                                                                            {4'b0010, 4'b0000, 4'b0000, 4'b0010, 4'b0100, 4'b0010, 4'b0010, 4'b1110, 4'b1110, 4'b0010, 4'b0010, 4'b0100, 4'b0010, 4'b1100, 4'b0100, 4'b0010, 4'b0000, 4'b1110, 4'b0000, 4'b0100, 4'b0100, 4'b1100, 4'b0010, 4'b0000, 4'b0010, 4'b0010, 4'b0010, 4'b0100, 4'b0010, 4'b0000, 4'b1110, 4'b0010},
                                                                                            {4'b0000, 4'b1110, 4'b1110, 4'b0100, 4'b0010, 4'b0100, 4'b0000, 4'b1100, 4'b1100, 4'b0000, 4'b0100, 4'b0010, 4'b0100, 4'b1110, 4'b0010, 4'b0100, 4'b1110, 4'b0000, 4'b1110, 4'b0010, 4'b0010, 4'b1110, 4'b0000, 4'b0010, 4'b0100, 4'b0000, 4'b0000, 4'b0010, 4'b0000, 4'b0010, 4'b0000, 4'b0000},
                                                                                            {4'b1110, 4'b0000, 4'b0000, 4'b1110, 4'b0000, 4'b1110, 4'b1110, 4'b0010, 4'b0010, 4'b1110, 4'b1110, 4'b0000, 4'b1110, 4'b0000, 4'b0000, 4'b1110, 4'b0100, 4'b0010, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0010, 4'b0000, 4'b1110, 4'b0010, 4'b1110, 4'b0000, 4'b0010, 4'b0000, 4'b0010, 4'b1110},
                                                                                            {4'b1100, 4'b1110, 4'b1110, 4'b0000, 4'b1110, 4'b0000, 4'b1100, 4'b0000, 4'b0000, 4'b1100, 4'b0000, 4'b1110, 4'b0000, 4'b0010, 4'b1110, 4'b0000, 4'b0010, 4'b0100, 4'b1110, 4'b1110, 4'b1110, 4'b0010, 4'b0000, 4'b0010, 4'b0000, 4'b0000, 4'b1100, 4'b1110, 4'b0000, 4'b0010, 4'b0100, 4'b1100},
                                                                                            {4'b0010, 4'b0100, 4'b0100, 4'b1110, 4'b0000, 4'b1110, 4'b0010, 4'b0010, 4'b0010, 4'b0010, 4'b1110, 4'b0000, 4'b1110, 4'b0000, 4'b0000, 4'b1110, 4'b0000, 4'b1110, 4'b0100, 4'b0000, 4'b0000, 4'b0000, 4'b0010, 4'b1100, 4'b1110, 4'b1110, 4'b0010, 4'b0000, 4'b1110, 4'b0000, 4'b1110, 4'b0010},
                                                                                            {4'b0010, 4'b0000, 4'b0000, 4'b0010, 4'b0100, 4'b0010, 4'b0010, 4'b1110, 4'b1110, 4'b0010, 4'b0010, 4'b0100, 4'b0010, 4'b1100, 4'b0100, 4'b0010, 4'b0000, 4'b1110, 4'b0000, 4'b0100, 4'b0100, 4'b1100, 4'b0010, 4'b0000, 4'b0010, 4'b0010, 4'b0010, 4'b0100, 4'b0010, 4'b0000, 4'b1110, 4'b0010},
                                                                                            {4'b0010, 4'b0000, 4'b0000, 4'b0010, 4'b0100, 4'b0010, 4'b0010, 4'b1110, 4'b1110, 4'b0010, 4'b0010, 4'b0100, 4'b0010, 4'b1100, 4'b0100, 4'b0010, 4'b0000, 4'b1110, 4'b0000, 4'b0100, 4'b0100, 4'b1100, 4'b0010, 4'b0000, 4'b0010, 4'b0010, 4'b0010, 4'b0100, 4'b0010, 4'b0000, 4'b1110, 4'b0010},
                                                                                            {4'b1110, 4'b0000, 4'b0000, 4'b1110, 4'b1100, 4'b1110, 4'b1110, 4'b0010, 4'b0010, 4'b1110, 4'b1110, 4'b1100, 4'b1110, 4'b0100, 4'b1100, 4'b1110, 4'b0000, 4'b0010, 4'b0000, 4'b1100, 4'b1100, 4'b0100, 4'b1110, 4'b0000, 4'b1110, 4'b1110, 4'b1110, 4'b1100, 4'b1110, 4'b0000, 4'b0010, 4'b1110},
                                                                                            {4'b0000, 4'b0010, 4'b0010, 4'b0000, 4'b0010, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0010, 4'b0000, 4'b1110, 4'b0010, 4'b0000, 4'b0010, 4'b0000, 4'b0010, 4'b0010, 4'b0010, 4'b1110, 4'b0100, 4'b1110, 4'b0000, 4'b0000, 4'b0000, 4'b0010, 4'b0000, 4'b0010, 4'b0000, 4'b0000},
                                                                                            {4'b1110, 4'b1100, 4'b1100, 4'b0010, 4'b0000, 4'b0010, 4'b1110, 4'b1110, 4'b1110, 4'b1110, 4'b0010, 4'b0000, 4'b0010, 4'b0000, 4'b0000, 4'b0010, 4'b0000, 4'b0010, 4'b1100, 4'b0000, 4'b0000, 4'b0000, 4'b1110, 4'b0100, 4'b0010, 4'b0010, 4'b1110, 4'b0000, 4'b0010, 4'b0000, 4'b0010, 4'b1110},
                                                                                            {4'b0000, 4'b1110, 4'b1110, 4'b0100, 4'b0010, 4'b0100, 4'b0000, 4'b1100, 4'b1100, 4'b0000, 4'b0100, 4'b0010, 4'b0100, 4'b1110, 4'b0010, 4'b0100, 4'b1110, 4'b0000, 4'b1110, 4'b0010, 4'b0010, 4'b1110, 4'b0000, 4'b0010, 4'b0100, 4'b0000, 4'b0000, 4'b0010, 4'b0000, 4'b0010, 4'b0000, 4'b0000},
                                                                                            {4'b0000, 4'b1110, 4'b1110, 4'b0000, 4'b0010, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0010, 4'b0000, 4'b1110, 4'b0010, 4'b0000, 4'b0010, 4'b0000, 4'b1110, 4'b0010, 4'b0010, 4'b1110, 4'b0000, 4'b0010, 4'b0000, 4'b0100, 4'b0000, 4'b0010, 4'b0100, 4'b1110, 4'b0000, 4'b0000},
                                                                                            {4'b0100, 4'b0010, 4'b0010, 4'b0000, 4'b0010, 4'b0000, 4'b0100, 4'b0000, 4'b0000, 4'b0100, 4'b0000, 4'b0010, 4'b0000, 4'b1110, 4'b0010, 4'b0000, 4'b1110, 4'b1100, 4'b0010, 4'b0010, 4'b0010, 4'b1110, 4'b0000, 4'b1110, 4'b0000, 4'b0000, 4'b0100, 4'b0010, 4'b0000, 4'b1110, 4'b1100, 4'b0100},
                                                                                            {4'b0010, 4'b0000, 4'b0000, 4'b0010, 4'b0100, 4'b0010, 4'b0010, 4'b1110, 4'b1110, 4'b0010, 4'b0010, 4'b0100, 4'b0010, 4'b1100, 4'b0100, 4'b0010, 4'b0000, 4'b1110, 4'b0000, 4'b0100, 4'b0100, 4'b1100, 4'b0010, 4'b0000, 4'b0010, 4'b0010, 4'b0010, 4'b0100, 4'b0010, 4'b0000, 4'b1110, 4'b0010},
                                                                                            {4'b0000, 4'b1110, 4'b1110, 4'b0000, 4'b0010, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0010, 4'b0000, 4'b1110, 4'b0010, 4'b0000, 4'b0010, 4'b0000, 4'b1110, 4'b0010, 4'b0010, 4'b1110, 4'b0000, 4'b0010, 4'b0000, 4'b0100, 4'b0000, 4'b0010, 4'b0100, 4'b1110, 4'b0000, 4'b0000},
                                                                                            {4'b1110, 4'b0000, 4'b0000, 4'b0010, 4'b0000, 4'b0010, 4'b1110, 4'b1110, 4'b1110, 4'b1110, 4'b0010, 4'b0000, 4'b0010, 4'b0000, 4'b0000, 4'b0010, 4'b0000, 4'b0010, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0010, 4'b0000, 4'b0010, 4'b1110, 4'b1110, 4'b0000, 4'b1110, 4'b0100, 4'b0010, 4'b1110},
                                                                                            {4'b1100, 4'b1110, 4'b1110, 4'b0000, 4'b1110, 4'b0000, 4'b1100, 4'b0000, 4'b0000, 4'b1100, 4'b0000, 4'b1110, 4'b0000, 4'b0010, 4'b1110, 4'b0000, 4'b0010, 4'b0100, 4'b1110, 4'b1110, 4'b1110, 4'b0010, 4'b0000, 4'b0010, 4'b0000, 4'b0000, 4'b1100, 4'b1110, 4'b0000, 4'b0010, 4'b0100, 4'b1100},
                                                                                            {4'b0100, 4'b0010, 4'b0010, 4'b0000, 4'b0010, 4'b0000, 4'b0100, 4'b0000, 4'b0000, 4'b0100, 4'b0000, 4'b0010, 4'b0000, 4'b1110, 4'b0010, 4'b0000, 4'b1110, 4'b1100, 4'b0010, 4'b0010, 4'b0010, 4'b1110, 4'b0000, 4'b1110, 4'b0000, 4'b0000, 4'b0100, 4'b0010, 4'b0000, 4'b1110, 4'b1100, 4'b0100}};



endpackage


`endif